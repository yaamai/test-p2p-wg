module chord

fn test_hoge() {
}
